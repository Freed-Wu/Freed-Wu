%FILE%
%HERE%
.end
