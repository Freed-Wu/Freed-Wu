module {{ expand('%:t:r') }};
  {% here %}
endmodule
